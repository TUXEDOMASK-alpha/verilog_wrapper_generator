module system_top (

);

    cpu cpu_inst (

    );

    memory mem_inst (

    );

endmodule